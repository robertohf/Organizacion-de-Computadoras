module DataMemory();
endmodule